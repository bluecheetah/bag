

module PYTEST(
    input  wire VDD,
    input  wire VSS,
    input  wire [3:0] vin,
    output wire vout
);

endmodule
