

module PYTEST(
    input  wire VDD,
    input  wire VSS,
    input  wire vin,
    output wire [3:0] mid,
    output wire vout
);

endmodule
